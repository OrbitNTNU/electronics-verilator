//add and substract
